<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>69.8879,-35.9607,119.894,-61.7513</PageViewport>
<gate>
<ID>2</ID>
<type>AE_DFF_LOW</type>
<position>86.5,-33</position>
<input>
<ID>IN_0</ID>4 </input>
<output>
<ID>OUTINV_0</ID>2 </output>
<output>
<ID>OUT_0</ID>1 </output>
<input>
<ID>clock</ID>3 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>79,-31</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>6</ID>
<type>GA_LED</type>
<position>93,-31</position>
<input>
<ID>N_in0</ID>1 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>7</ID>
<type>GA_LED</type>
<position>93,-34</position>
<input>
<ID>N_in0</ID>2 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>79,-34</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>9</ID>
<type>AA_TOGGLE</type>
<position>74,-43</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>74,-49</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>14</ID>
<type>BA_NAND2</type>
<position>88,-45</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>15</ID>
<type>BA_NAND2</type>
<position>99,-46</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>5 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>16</ID>
<type>BA_NAND2</type>
<position>99,-52</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>17</ID>
<type>BA_NAND2</type>
<position>88,-53</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>18</ID>
<type>GA_LED</type>
<position>106,-46</position>
<input>
<ID>N_in0</ID>6 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>GA_LED</type>
<position>106,-52</position>
<input>
<ID>N_in0</ID>5 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>21</ID>
<type>AE_SMALL_INVERTER</type>
<position>82,-54</position>
<input>
<ID>IN_0</ID>8 </input>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>89.5,-31,92,-31</points>
<connection>
<GID>6</GID>
<name>N_in0</name></connection>
<intersection>89.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>89.5,-31,89.5,-31</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>-31 1</intersection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>89.5,-34,92,-34</points>
<connection>
<GID>2</GID>
<name>OUTINV_0</name></connection>
<connection>
<GID>7</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>81,-34,83.5,-34</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<connection>
<GID>2</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>81,-31,83.5,-31</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>95,-48.5,104,-48.5</points>
<intersection>95 3</intersection>
<intersection>104 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>95,-48.5,95,-47</points>
<intersection>-48.5 1</intersection>
<intersection>-47 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>95,-47,96,-47</points>
<connection>
<GID>15</GID>
<name>IN_1</name></connection>
<intersection>95 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>104,-52,104,-48.5</points>
<intersection>-52 7</intersection>
<intersection>-48.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>102,-52,105,-52</points>
<connection>
<GID>19</GID>
<name>N_in0</name></connection>
<connection>
<GID>16</GID>
<name>OUT</name></connection>
<intersection>104 5</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94,-49.5,103,-49.5</points>
<intersection>94 3</intersection>
<intersection>103 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>94,-51,94,-49.5</points>
<intersection>-51 4</intersection>
<intersection>-49.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>94,-51,96,-51</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>94 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>103,-49.5,103,-46</points>
<intersection>-49.5 1</intersection>
<intersection>-46 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>102,-46,105,-46</points>
<connection>
<GID>18</GID>
<name>N_in0</name></connection>
<connection>
<GID>15</GID>
<name>OUT</name></connection>
<intersection>103 5</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>84,-54,85,-54</points>
<connection>
<GID>21</GID>
<name>OUT_0</name></connection>
<connection>
<GID>17</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79,-54,79,-43</points>
<intersection>-54 2</intersection>
<intersection>-44 3</intersection>
<intersection>-43 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76,-43,79,-43</points>
<connection>
<GID>9</GID>
<name>OUT_0</name></connection>
<intersection>79 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>79,-54,80,-54</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>79 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>79,-44,85,-44</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>79 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81,-52,81,-46</points>
<intersection>-52 3</intersection>
<intersection>-49 1</intersection>
<intersection>-46 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76,-49,81,-49</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>81,-46,85,-46</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>81,-52,85,-52</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<intersection>81 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>91,-45,96,-45</points>
<connection>
<GID>14</GID>
<name>OUT</name></connection>
<connection>
<GID>15</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>91,-53,96,-53</points>
<connection>
<GID>17</GID>
<name>OUT</name></connection>
<connection>
<GID>16</GID>
<name>IN_1</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,177.8,-91.7</PageViewport></page 1>
<page 2>
<PageViewport>0,0,177.8,-91.7</PageViewport></page 2>
<page 3>
<PageViewport>0,0,177.8,-91.7</PageViewport></page 3>
<page 4>
<PageViewport>0,0,177.8,-91.7</PageViewport></page 4>
<page 5>
<PageViewport>0,0,177.8,-91.7</PageViewport></page 5>
<page 6>
<PageViewport>0,0,177.8,-91.7</PageViewport></page 6>
<page 7>
<PageViewport>0,0,177.8,-91.7</PageViewport></page 7>
<page 8>
<PageViewport>0,0,177.8,-91.7</PageViewport></page 8>
<page 9>
<PageViewport>0,0,177.8,-91.7</PageViewport></page 9></circuit>